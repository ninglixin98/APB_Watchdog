`ifndef RKV_WATCHDOG_CONFIG_SVH
`define RKV_WATCHDOG_CONFIG_SVH

`include "rkv_watchdog_config.sv"

`endif//RKV_WATCHDOG_CONFIG_SVH

